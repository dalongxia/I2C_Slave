module i2c_slave_top(
	input	clk,
	input	rst_n,
	input	scl,
	inout	sda,
	output	dav,
	output	dout

);


endmodule
